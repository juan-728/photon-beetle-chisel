module Photon(
  input        clock,
  input        reset,
  input  [7:0] io_state_0_0,
  input  [7:0] io_state_0_1,
  input  [7:0] io_state_0_2,
  input  [7:0] io_state_0_3,
  input  [7:0] io_state_0_4,
  input  [7:0] io_state_0_5,
  input  [7:0] io_state_0_6,
  input  [7:0] io_state_0_7,
  input  [7:0] io_state_1_0,
  input  [7:0] io_state_1_1,
  input  [7:0] io_state_1_2,
  input  [7:0] io_state_1_3,
  input  [7:0] io_state_1_4,
  input  [7:0] io_state_1_5,
  input  [7:0] io_state_1_6,
  input  [7:0] io_state_1_7,
  input  [7:0] io_state_2_0,
  input  [7:0] io_state_2_1,
  input  [7:0] io_state_2_2,
  input  [7:0] io_state_2_3,
  input  [7:0] io_state_2_4,
  input  [7:0] io_state_2_5,
  input  [7:0] io_state_2_6,
  input  [7:0] io_state_2_7,
  input  [7:0] io_state_3_0,
  input  [7:0] io_state_3_1,
  input  [7:0] io_state_3_2,
  input  [7:0] io_state_3_3,
  input  [7:0] io_state_3_4,
  input  [7:0] io_state_3_5,
  input  [7:0] io_state_3_6,
  input  [7:0] io_state_3_7,
  input  [7:0] io_state_4_0,
  input  [7:0] io_state_4_1,
  input  [7:0] io_state_4_2,
  input  [7:0] io_state_4_3,
  input  [7:0] io_state_4_4,
  input  [7:0] io_state_4_5,
  input  [7:0] io_state_4_6,
  input  [7:0] io_state_4_7,
  input  [7:0] io_state_5_0,
  input  [7:0] io_state_5_1,
  input  [7:0] io_state_5_2,
  input  [7:0] io_state_5_3,
  input  [7:0] io_state_5_4,
  input  [7:0] io_state_5_5,
  input  [7:0] io_state_5_6,
  input  [7:0] io_state_5_7,
  input  [7:0] io_state_6_0,
  input  [7:0] io_state_6_1,
  input  [7:0] io_state_6_2,
  input  [7:0] io_state_6_3,
  input  [7:0] io_state_6_4,
  input  [7:0] io_state_6_5,
  input  [7:0] io_state_6_6,
  input  [7:0] io_state_6_7,
  input  [7:0] io_state_7_0,
  input  [7:0] io_state_7_1,
  input  [7:0] io_state_7_2,
  input  [7:0] io_state_7_3,
  input  [7:0] io_state_7_4,
  input  [7:0] io_state_7_5,
  input  [7:0] io_state_7_6,
  input  [7:0] io_state_7_7
);
endmodule
