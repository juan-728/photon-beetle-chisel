module Photon_Beetle_HASH(
  input         clock,
  input         reset,
  input  [3:0]  io_state_0_0,
  input  [3:0]  io_state_0_1,
  input  [3:0]  io_state_0_2,
  input  [3:0]  io_state_0_3,
  input  [3:0]  io_state_0_4,
  input  [3:0]  io_state_0_5,
  input  [3:0]  io_state_0_6,
  input  [3:0]  io_state_0_7,
  input  [3:0]  io_state_1_0,
  input  [3:0]  io_state_1_1,
  input  [3:0]  io_state_1_2,
  input  [3:0]  io_state_1_3,
  input  [3:0]  io_state_1_4,
  input  [3:0]  io_state_1_5,
  input  [3:0]  io_state_1_6,
  input  [3:0]  io_state_1_7,
  input  [3:0]  io_state_2_0,
  input  [3:0]  io_state_2_1,
  input  [3:0]  io_state_2_2,
  input  [3:0]  io_state_2_3,
  input  [3:0]  io_state_2_4,
  input  [3:0]  io_state_2_5,
  input  [3:0]  io_state_2_6,
  input  [3:0]  io_state_2_7,
  input  [3:0]  io_state_3_0,
  input  [3:0]  io_state_3_1,
  input  [3:0]  io_state_3_2,
  input  [3:0]  io_state_3_3,
  input  [3:0]  io_state_3_4,
  input  [3:0]  io_state_3_5,
  input  [3:0]  io_state_3_6,
  input  [3:0]  io_state_3_7,
  input  [3:0]  io_state_4_0,
  input  [3:0]  io_state_4_1,
  input  [3:0]  io_state_4_2,
  input  [3:0]  io_state_4_3,
  input  [3:0]  io_state_4_4,
  input  [3:0]  io_state_4_5,
  input  [3:0]  io_state_4_6,
  input  [3:0]  io_state_4_7,
  input  [3:0]  io_state_5_0,
  input  [3:0]  io_state_5_1,
  input  [3:0]  io_state_5_2,
  input  [3:0]  io_state_5_3,
  input  [3:0]  io_state_5_4,
  input  [3:0]  io_state_5_5,
  input  [3:0]  io_state_5_6,
  input  [3:0]  io_state_5_7,
  input  [3:0]  io_state_6_0,
  input  [3:0]  io_state_6_1,
  input  [3:0]  io_state_6_2,
  input  [3:0]  io_state_6_3,
  input  [3:0]  io_state_6_4,
  input  [3:0]  io_state_6_5,
  input  [3:0]  io_state_6_6,
  input  [3:0]  io_state_6_7,
  input  [3:0]  io_state_7_0,
  input  [3:0]  io_state_7_1,
  input  [3:0]  io_state_7_2,
  input  [3:0]  io_state_7_3,
  input  [3:0]  io_state_7_4,
  input  [3:0]  io_state_7_5,
  input  [3:0]  io_state_7_6,
  input  [3:0]  io_state_7_7,
  input         io_condition,
  input  [7:0]  io_option1,
  input  [7:0]  io_option2,
  input  [7:0]  io_out_0,
  input  [7:0]  io_out_1,
  input  [7:0]  io_out_2,
  input  [7:0]  io_out_3,
  input  [7:0]  io_in,
  input  [7:0]  io_in_left_0,
  input  [7:0]  io_in_left_1,
  input  [7:0]  io_in_left_2,
  input  [7:0]  io_in_left_3,
  input  [7:0]  io_in_right_0,
  input  [7:0]  io_in_right_1,
  input  [7:0]  io_in_right_2,
  input  [7:0]  io_in_right_3,
  input  [31:0] io_iolen_inbytes,
  input  [63:0] io_inlen,
  input  [3:0]  io_State_inout_0,
  input  [3:0]  io_State_inout_1,
  input  [3:0]  io_State_inout_2,
  input  [3:0]  io_State_inout_3,
  input  [3:0]  io_State_inout_4,
  input  [3:0]  io_State_inout_5,
  input  [3:0]  io_State_inout_6,
  input  [3:0]  io_State_inout_7,
  input  [3:0]  io_State_inout_8,
  input  [3:0]  io_State_inout_9,
  input  [3:0]  io_State_inout_10,
  input  [3:0]  io_State_inout_11,
  input  [3:0]  io_State_inout_12,
  input  [3:0]  io_State_inout_13,
  input  [3:0]  io_State_inout_14,
  input  [3:0]  io_State_inout_15,
  input  [3:0]  io_State_inout_16,
  input  [3:0]  io_State_inout_17,
  input  [3:0]  io_State_inout_18,
  input  [3:0]  io_State_inout_19,
  input  [3:0]  io_State_inout_20,
  input  [3:0]  io_State_inout_21,
  input  [3:0]  io_State_inout_22,
  input  [3:0]  io_State_inout_23,
  input  [3:0]  io_State_inout_24,
  input  [3:0]  io_State_inout_25,
  input  [3:0]  io_State_inout_26,
  input  [3:0]  io_State_inout_27,
  input  [3:0]  io_State_inout_28,
  input  [3:0]  io_State_inout_29,
  input  [3:0]  io_State_inout_30,
  input  [3:0]  io_State_inout_31,
  input  [3:0]  io_State_inout_32,
  input  [3:0]  io_State_inout_33,
  input  [3:0]  io_State_inout_34,
  input  [3:0]  io_State_inout_35,
  input  [3:0]  io_State_inout_36,
  input  [3:0]  io_State_inout_37,
  input  [3:0]  io_State_inout_38,
  input  [3:0]  io_State_inout_39,
  input  [3:0]  io_State_inout_40,
  input  [3:0]  io_State_inout_41,
  input  [3:0]  io_State_inout_42,
  input  [3:0]  io_State_inout_43,
  input  [3:0]  io_State_inout_44,
  input  [3:0]  io_State_inout_45,
  input  [3:0]  io_State_inout_46,
  input  [3:0]  io_State_inout_47,
  input  [3:0]  io_State_inout_48,
  input  [3:0]  io_State_inout_49,
  input  [3:0]  io_State_inout_50,
  input  [3:0]  io_State_inout_51,
  input  [3:0]  io_State_inout_52,
  input  [3:0]  io_State_inout_53,
  input  [3:0]  io_State_inout_54,
  input  [3:0]  io_State_inout_55,
  input  [3:0]  io_State_inout_56,
  input  [3:0]  io_State_inout_57,
  input  [3:0]  io_State_inout_58,
  input  [3:0]  io_State_inout_59,
  input  [3:0]  io_State_inout_60,
  input  [3:0]  io_State_inout_61,
  input  [3:0]  io_State_inout_62,
  input  [3:0]  io_State_inout_63,
  input  [7:0]  io_Constant,
  input  [7:0]  io_Data_in_0,
  input  [7:0]  io_Data_in_1,
  input  [7:0]  io_Data_in_2,
  input  [7:0]  io_Data_in_3,
  input  [63:0] io_Dlen_inbytes,
  input  [7:0]  io_State,
  input  [7:0]  io_Tag_out_0,
  input  [7:0]  io_Tag_out_1,
  input  [7:0]  io_Tag_out_2,
  input  [7:0]  io_Tag_out_3,
  input  [7:0]  io_Tag_out_4,
  input  [7:0]  io_Tag_out_5,
  input  [7:0]  io_Tag_out_6,
  input  [7:0]  io_Tag_out_7,
  input  [7:0]  io_Tag_out_8,
  input  [7:0]  io_Tag_out_9,
  input  [7:0]  io_Tag_out_10,
  input  [7:0]  io_Tag_out_11,
  input  [7:0]  io_Tag_out_12,
  input  [7:0]  io_Tag_out_13,
  input  [7:0]  io_Tag_out_14,
  input  [7:0]  io_Tag_out_15,
  input  [3:0]  io_state_in_0,
  input  [3:0]  io_state_in_1,
  input  [3:0]  io_state_in_2,
  input  [3:0]  io_state_in_3,
  input  [3:0]  io_state_in_4,
  input  [3:0]  io_state_in_5,
  input  [3:0]  io_state_in_6,
  input  [3:0]  io_state_in_7,
  input  [3:0]  io_state_in_8,
  input  [3:0]  io_state_in_9,
  input  [3:0]  io_state_in_10,
  input  [3:0]  io_state_in_11,
  input  [3:0]  io_state_in_12,
  input  [3:0]  io_state_in_13,
  input  [3:0]  io_state_in_14,
  input  [3:0]  io_state_in_15,
  input  [3:0]  io_state_in_16,
  input  [3:0]  io_state_in_17,
  input  [3:0]  io_state_in_18,
  input  [3:0]  io_state_in_19,
  input  [3:0]  io_state_in_20,
  input  [3:0]  io_state_in_21,
  input  [3:0]  io_state_in_22,
  input  [3:0]  io_state_in_23,
  input  [3:0]  io_state_in_24,
  input  [3:0]  io_state_in_25,
  input  [3:0]  io_state_in_26,
  input  [3:0]  io_state_in_27,
  input  [3:0]  io_state_in_28,
  input  [3:0]  io_state_in_29,
  input  [3:0]  io_state_in_30,
  input  [3:0]  io_state_in_31,
  input  [3:0]  io_state_in_32,
  input  [3:0]  io_state_in_33,
  input  [3:0]  io_state_in_34,
  input  [3:0]  io_state_in_35,
  input  [3:0]  io_state_in_36,
  input  [3:0]  io_state_in_37,
  input  [3:0]  io_state_in_38,
  input  [3:0]  io_state_in_39,
  input  [3:0]  io_state_in_40,
  input  [3:0]  io_state_in_41,
  input  [3:0]  io_state_in_42,
  input  [3:0]  io_state_in_43,
  input  [3:0]  io_state_in_44,
  input  [3:0]  io_state_in_45,
  input  [3:0]  io_state_in_46,
  input  [3:0]  io_state_in_47,
  input  [3:0]  io_state_in_48,
  input  [3:0]  io_state_in_49,
  input  [3:0]  io_state_in_50,
  input  [3:0]  io_state_in_51,
  input  [3:0]  io_state_in_52,
  input  [3:0]  io_state_in_53,
  input  [3:0]  io_state_in_54,
  input  [3:0]  io_state_in_55,
  input  [3:0]  io_state_in_56,
  input  [3:0]  io_state_in_57,
  input  [3:0]  io_state_in_58,
  input  [3:0]  io_state_in_59,
  input  [3:0]  io_state_in_60,
  input  [3:0]  io_state_in_61,
  input  [3:0]  io_state_in_62,
  input  [3:0]  io_state_in_63,
  input  [3:0]  io_state_out_0,
  input  [3:0]  io_state_out_1,
  input  [3:0]  io_state_out_2,
  input  [3:0]  io_state_out_3,
  input  [3:0]  io_state_out_4,
  input  [3:0]  io_state_out_5,
  input  [3:0]  io_state_out_6,
  input  [3:0]  io_state_out_7,
  input  [3:0]  io_state_out_8,
  input  [3:0]  io_state_out_9,
  input  [3:0]  io_state_out_10,
  input  [3:0]  io_state_out_11,
  input  [3:0]  io_state_out_12,
  input  [3:0]  io_state_out_13,
  input  [3:0]  io_state_out_14,
  input  [3:0]  io_state_out_15,
  input  [3:0]  io_state_out_16,
  input  [3:0]  io_state_out_17,
  input  [3:0]  io_state_out_18,
  input  [3:0]  io_state_out_19,
  input  [3:0]  io_state_out_20,
  input  [3:0]  io_state_out_21,
  input  [3:0]  io_state_out_22,
  input  [3:0]  io_state_out_23,
  input  [3:0]  io_state_out_24,
  input  [3:0]  io_state_out_25,
  input  [3:0]  io_state_out_26,
  input  [3:0]  io_state_out_27,
  input  [3:0]  io_state_out_28,
  input  [3:0]  io_state_out_29,
  input  [3:0]  io_state_out_30,
  input  [3:0]  io_state_out_31,
  input  [3:0]  io_state_out_32,
  input  [3:0]  io_state_out_33,
  input  [3:0]  io_state_out_34,
  input  [3:0]  io_state_out_35,
  input  [3:0]  io_state_out_36,
  input  [3:0]  io_state_out_37,
  input  [3:0]  io_state_out_38,
  input  [3:0]  io_state_out_39,
  input  [3:0]  io_state_out_40,
  input  [3:0]  io_state_out_41,
  input  [3:0]  io_state_out_42,
  input  [3:0]  io_state_out_43,
  input  [3:0]  io_state_out_44,
  input  [3:0]  io_state_out_45,
  input  [3:0]  io_state_out_46,
  input  [3:0]  io_state_out_47,
  input  [3:0]  io_state_out_48,
  input  [3:0]  io_state_out_49,
  input  [3:0]  io_state_out_50,
  input  [3:0]  io_state_out_51,
  input  [3:0]  io_state_out_52,
  input  [3:0]  io_state_out_53,
  input  [3:0]  io_state_out_54,
  input  [3:0]  io_state_out_55,
  input  [3:0]  io_state_out_56,
  input  [3:0]  io_state_out_57,
  input  [3:0]  io_state_out_58,
  input  [3:0]  io_state_out_59,
  input  [3:0]  io_state_out_60,
  input  [3:0]  io_state_out_61,
  input  [3:0]  io_state_out_62,
  input  [3:0]  io_state_out_63,
  input  [31:0] io_round
);
endmodule
